magic
tech scmos
timestamp 1668616580
<< metal1 >>
rect -77 77 -15 81
rect -10 77 111 81
rect 116 77 489 81
rect 494 77 867 81
rect 872 77 2038 81
rect -77 66 237 70
rect 242 66 615 70
rect 620 66 741 70
rect 746 66 1371 70
rect 1376 66 2035 70
rect -77 55 363 59
rect 368 55 1119 59
rect 1124 55 1245 59
rect 1250 55 1623 59
rect 1628 55 2038 59
rect -77 44 993 48
rect 998 44 1497 48
rect 1502 44 1749 48
rect 1754 44 1875 48
rect 1880 44 2038 48
rect -77 33 -29 37
rect -24 33 223 37
rect 228 33 349 37
rect 354 33 979 37
rect 984 33 2036 37
rect -77 22 97 26
rect 102 22 601 26
rect 606 22 1105 26
rect 1110 22 1483 26
rect 1488 22 2039 26
rect -77 11 475 15
rect 480 11 727 15
rect 732 11 1231 15
rect 1236 11 1735 15
rect 1740 11 2038 15
rect -77 0 853 4
rect 858 0 1357 4
rect 1362 0 1609 4
rect 1614 0 1861 4
rect 1866 0 2038 4
rect 1883 -52 1884 -51
rect -77 -56 -5 -52
rect 48 -56 122 -52
rect 174 -56 248 -52
rect 300 -56 374 -52
rect 425 -56 499 -52
rect 550 -56 625 -52
rect 678 -56 753 -52
rect 804 -56 879 -52
rect 931 -56 1006 -52
rect 1056 -56 1131 -52
rect 1182 -56 1257 -52
rect 1309 -56 1384 -52
rect 1435 -56 1510 -52
rect 1561 -56 1636 -52
rect 1687 -56 1762 -52
rect 1813 -55 1888 -52
rect 1813 -56 1883 -55
rect -10 -81 -6 -77
rect 116 -81 121 -77
rect 242 -81 246 -77
rect 368 -81 372 -77
rect 494 -81 498 -77
rect 620 -81 624 -77
rect 746 -81 750 -77
rect 871 -81 876 -77
rect 998 -81 1002 -77
rect 1124 -81 1128 -77
rect 1250 -81 1254 -77
rect 1376 -81 1380 -77
rect 1502 -81 1506 -77
rect 1628 -81 1632 -77
rect 1754 -81 1758 -77
rect 1880 -80 1884 -76
rect -24 -88 -6 -84
rect 49 -89 65 -85
rect 102 -88 121 -84
rect 176 -89 191 -85
rect 228 -88 246 -84
rect 302 -89 317 -85
rect 354 -88 372 -84
rect 428 -89 443 -85
rect 480 -88 498 -84
rect 554 -89 569 -85
rect 606 -88 624 -84
rect 680 -89 695 -85
rect 732 -88 750 -84
rect 806 -89 821 -85
rect 858 -88 876 -84
rect 932 -89 947 -85
rect 984 -88 1002 -84
rect 1058 -89 1073 -85
rect 1110 -88 1128 -84
rect 1184 -89 1199 -85
rect 1236 -88 1254 -84
rect 1310 -89 1325 -85
rect 1362 -88 1380 -84
rect 1436 -89 1451 -85
rect 1488 -88 1506 -84
rect 1562 -89 1577 -85
rect 1614 -88 1632 -84
rect 1688 -89 1703 -85
rect 1740 -88 1758 -84
rect 1814 -89 1829 -85
rect 1866 -87 1884 -83
rect 1940 -88 1955 -84
rect -77 -110 -6 -106
rect 61 -378 65 -89
rect -676 -382 65 -378
rect -676 -2388 -672 -382
rect 187 -449 191 -89
rect -612 -453 191 -449
rect -612 -637 -608 -453
rect 313 -473 317 -89
rect 439 -364 443 -89
rect -585 -477 317 -473
rect 388 -368 443 -364
rect -585 -616 -581 -477
rect 342 -593 353 -589
rect -585 -620 -545 -616
rect -612 -641 -543 -637
rect -635 -797 -543 -793
rect 340 -1361 344 -703
rect 91 -1365 344 -1361
rect -470 -1844 80 -1840
rect -470 -2359 -466 -1844
rect 91 -1873 95 -1365
rect -438 -1877 95 -1873
rect 112 -1381 379 -1377
rect -438 -2247 -434 -1877
rect 112 -1916 116 -1381
rect 388 -1450 392 -368
rect 439 -632 443 -379
rect 435 -636 443 -632
rect 435 -1006 439 -636
rect 565 -650 569 -89
rect 691 -193 695 -89
rect 817 -219 821 -89
rect 700 -223 821 -219
rect 700 -402 704 -223
rect 943 -229 947 -89
rect 731 -233 947 -229
rect 731 -381 735 -233
rect 970 -316 1002 -312
rect 731 -385 768 -381
rect 700 -406 766 -402
rect 969 -470 982 -466
rect 1069 -572 1073 -89
rect 1195 -131 1199 -89
rect 1127 -135 1199 -131
rect 1321 -219 1325 -89
rect 1189 -223 1325 -219
rect 1189 -403 1193 -223
rect 1447 -229 1451 -89
rect 1224 -233 1451 -229
rect 1224 -382 1228 -233
rect 1460 -317 1499 -313
rect 1224 -386 1260 -382
rect 1189 -407 1257 -403
rect 1462 -471 1473 -467
rect 1069 -576 1555 -572
rect 646 -618 1492 -614
rect 445 -654 569 -650
rect 445 -850 449 -654
rect 1488 -802 1492 -618
rect 1374 -806 1492 -802
rect 462 -833 506 -829
rect 445 -854 506 -850
rect 1391 -920 1404 -916
rect 435 -1010 508 -1006
rect 1400 -1173 1404 -920
rect 1429 -1154 1534 -1150
rect 1551 -1166 1555 -576
rect 1573 -1068 1577 -89
rect 1699 -219 1703 -89
rect 1688 -223 1703 -219
rect 1688 -403 1692 -223
rect 1825 -229 1829 -89
rect 1951 -126 1955 -88
rect 1951 -130 4016 -126
rect 1724 -233 1829 -229
rect 1724 -382 1728 -233
rect 1973 -317 2025 -313
rect 1724 -386 1770 -382
rect 1688 -407 1769 -403
rect 1973 -471 1992 -467
rect 3377 -1024 3405 -1020
rect 1998 -1051 2494 -1047
rect 1573 -1072 2497 -1068
rect 3377 -1138 3405 -1134
rect 1551 -1170 2348 -1166
rect 1277 -1196 1505 -1192
rect 186 -1454 392 -1450
rect 186 -1596 190 -1454
rect 1094 -1569 1098 -1382
rect 1277 -1529 1281 -1196
rect 1309 -1209 1472 -1205
rect 1309 -1373 1313 -1209
rect 2228 -1329 2232 -1183
rect 1337 -1356 1344 -1352
rect 1309 -1377 1344 -1373
rect 1277 -1533 1343 -1529
rect 1092 -1573 1098 -1569
rect 1610 -1586 1675 -1582
rect 186 -1600 208 -1596
rect 180 -1621 210 -1617
rect 1079 -1687 1380 -1683
rect 167 -1777 210 -1773
rect 128 -1844 542 -1840
rect -393 -1920 116 -1916
rect -393 -2070 -389 -1920
rect 538 -2043 542 -1844
rect 522 -2047 542 -2043
rect -393 -2074 -361 -2070
rect -414 -2095 -361 -2091
rect 673 -2104 677 -1864
rect 1358 -2012 1362 -1897
rect 1376 -1917 1380 -1687
rect 1610 -1780 1614 -1586
rect 2226 -1702 2230 -1439
rect 2161 -1706 2230 -1702
rect 1673 -1831 1699 -1827
rect 2161 -1876 2165 -1706
rect 2344 -1713 2348 -1170
rect 2483 -1228 2496 -1224
rect 2401 -1653 3082 -1649
rect 2172 -1717 2348 -1713
rect 2172 -1855 2176 -1717
rect 3078 -1832 3082 -1653
rect 2172 -1859 2195 -1855
rect 2161 -1880 2194 -1876
rect 1437 -1900 1474 -1896
rect 1376 -1921 1473 -1917
rect 3075 -1946 3103 -1942
rect 1675 -1985 1696 -1981
rect 1692 -2012 1696 -1985
rect 1358 -2016 1696 -2012
rect 2151 -2036 2195 -2032
rect 405 -2108 677 -2104
rect 514 -2161 546 -2157
rect -438 -2251 -358 -2247
rect -1376 -2392 -672 -2388
rect -1376 -2530 -1372 -2392
rect -466 -2507 -441 -2503
rect -1376 -2534 -1348 -2530
rect -1383 -2555 -1346 -2551
rect 4012 -2557 4016 -130
rect -470 -2621 -436 -2617
rect -1392 -2711 -1349 -2707
<< m2contact >>
rect -15 76 -10 81
rect 111 76 116 81
rect 489 76 494 81
rect 867 76 872 81
rect 237 65 242 70
rect 615 65 620 70
rect 741 65 746 70
rect 1371 65 1376 70
rect 363 54 368 59
rect 1119 54 1124 59
rect 1245 54 1250 59
rect 1623 54 1628 59
rect 993 43 998 48
rect 1497 43 1502 48
rect 1749 43 1754 48
rect 1875 43 1880 48
rect -29 32 -24 37
rect 223 32 228 37
rect 349 32 354 37
rect 979 32 984 37
rect 97 21 102 26
rect 601 21 606 26
rect 1105 21 1110 26
rect 1483 21 1488 26
rect 475 10 480 15
rect 727 10 732 15
rect 1231 10 1236 15
rect 1735 10 1740 15
rect 853 -1 858 4
rect 1357 -1 1362 4
rect 1609 -1 1614 4
rect 1861 -1 1866 4
rect -15 -81 -10 -76
rect 111 -81 116 -76
rect 237 -81 242 -76
rect 363 -81 368 -76
rect 489 -81 494 -76
rect 615 -81 620 -76
rect 741 -81 746 -76
rect 866 -81 871 -76
rect 993 -81 998 -76
rect 1119 -81 1124 -76
rect 1245 -81 1250 -76
rect 1371 -81 1376 -76
rect 1497 -81 1502 -76
rect 1623 -81 1628 -76
rect 1749 -81 1754 -76
rect 1875 -80 1880 -75
rect -29 -88 -24 -83
rect 97 -88 102 -83
rect 223 -88 228 -83
rect 349 -88 354 -83
rect 475 -88 480 -83
rect 601 -88 606 -83
rect 727 -88 732 -83
rect 853 -88 858 -83
rect 979 -88 984 -83
rect 1105 -88 1110 -83
rect 1231 -88 1236 -83
rect 1357 -88 1362 -83
rect 1483 -88 1488 -83
rect 1609 -88 1614 -83
rect 1735 -88 1740 -83
rect 1861 -87 1866 -82
rect 46 -111 52 -106
rect 118 -111 124 -106
rect 173 -111 179 -106
rect 244 -111 250 -106
rect 300 -111 306 -106
rect 426 -111 432 -106
rect 496 -111 502 -106
rect 550 -111 556 -106
rect 353 -594 358 -589
rect -640 -797 -635 -792
rect 80 -1846 86 -1839
rect 379 -1382 384 -1377
rect 439 -379 444 -374
rect 622 -111 628 -106
rect 676 -111 682 -106
rect 748 -111 754 -106
rect 803 -111 809 -106
rect 690 -198 695 -193
rect 873 -111 879 -106
rect 928 -111 934 -106
rect 1000 -111 1006 -106
rect 1055 -111 1061 -106
rect 1002 -317 1007 -312
rect 982 -471 987 -466
rect 1125 -111 1131 -106
rect 1252 -111 1258 -106
rect 1308 -111 1314 -106
rect 1122 -136 1127 -131
rect 1379 -111 1385 -106
rect 1432 -111 1438 -106
rect 1504 -111 1510 -106
rect 1559 -111 1565 -106
rect 1499 -318 1504 -313
rect 1473 -472 1478 -467
rect 641 -618 646 -613
rect 457 -833 462 -828
rect 1421 -1154 1429 -1149
rect 1534 -1155 1541 -1150
rect 1630 -111 1636 -106
rect 1685 -111 1691 -106
rect 1757 -111 1763 -106
rect 1812 -111 1818 -106
rect 1881 -110 1887 -105
rect 2025 -318 2030 -313
rect 1992 -472 1997 -467
rect 3405 -1024 3410 -1019
rect 1993 -1051 1998 -1046
rect 1399 -1178 1404 -1173
rect 2228 -1183 2233 -1178
rect 1505 -1196 1510 -1191
rect 1093 -1382 1098 -1377
rect 1472 -1209 1477 -1204
rect 1332 -1356 1337 -1351
rect 175 -1621 180 -1616
rect 162 -1777 167 -1772
rect 122 -1846 128 -1840
rect 673 -1864 678 -1859
rect -419 -2095 -414 -2090
rect 400 -2108 405 -2103
rect 1357 -1897 1362 -1892
rect 2478 -1228 2483 -1223
rect 2395 -1653 2401 -1648
rect 1432 -1900 1437 -1895
rect 2146 -2036 2151 -2031
rect -471 -2364 -466 -2359
rect -1388 -2555 -1383 -2550
rect -1397 -2711 -1392 -2706
<< metal2 >>
rect -29 -83 -25 32
rect -15 -76 -11 76
rect 97 -83 101 21
rect 111 -76 115 76
rect 223 -83 227 32
rect 237 -76 241 65
rect 349 -83 353 32
rect 363 -76 367 54
rect 475 -83 479 10
rect 489 -76 493 76
rect 601 -83 605 21
rect 615 -76 619 65
rect 727 -83 731 10
rect 741 -76 745 65
rect 853 -83 857 -1
rect 867 -76 871 76
rect 979 -83 983 32
rect 993 -76 997 43
rect 1105 -83 1109 21
rect 1119 -76 1123 54
rect 1231 -83 1235 10
rect 1245 -76 1249 54
rect 1357 -83 1361 -1
rect 1371 -76 1375 65
rect 1483 -83 1487 21
rect 1497 -76 1501 43
rect 1609 -83 1613 -1
rect 1623 -76 1627 54
rect 1735 -83 1739 10
rect 1749 -76 1753 43
rect 1861 -82 1865 -1
rect 1875 -75 1879 43
rect 52 -110 118 -106
rect 179 -110 244 -106
rect 306 -110 375 -106
rect 432 -110 496 -106
rect 556 -110 622 -106
rect 682 -110 748 -106
rect 809 -110 873 -106
rect 934 -110 1000 -106
rect 1061 -110 1125 -106
rect 1187 -110 1252 -106
rect 1314 -110 1379 -106
rect 1438 -110 1504 -106
rect 1565 -110 1630 -106
rect 1691 -110 1757 -106
rect 1818 -110 1881 -106
rect 599 -198 690 -194
rect 599 -374 603 -198
rect 444 -378 603 -374
rect -640 -405 645 -401
rect -640 -792 -636 -405
rect -117 -489 619 -485
rect 354 -1130 358 -594
rect 641 -613 645 -405
rect 763 -489 852 -485
rect 983 -668 987 -471
rect 457 -672 987 -668
rect 1003 -667 1007 -317
rect 1122 -638 1126 -136
rect 1474 -589 1478 -472
rect 1500 -574 1504 -318
rect 1654 -493 1857 -489
rect 1500 -578 1529 -574
rect 1474 -593 1510 -589
rect 1122 -642 1477 -638
rect 1003 -671 1466 -667
rect 457 -828 461 -672
rect 329 -1134 358 -1130
rect 329 -1353 333 -1134
rect 68 -1357 333 -1353
rect 358 -1154 1421 -1150
rect 68 -1855 72 -1357
rect 358 -1423 362 -1154
rect 162 -1427 362 -1423
rect 371 -1178 1399 -1174
rect 162 -1772 166 -1427
rect 371 -1436 375 -1178
rect 1462 -1214 1466 -671
rect 1473 -1204 1477 -642
rect 1506 -1191 1510 -593
rect 1525 -1192 1529 -578
rect 1993 -1046 1997 -472
rect 2026 -512 2030 -318
rect 2534 -911 3410 -907
rect 1541 -1154 2232 -1150
rect 2228 -1178 2232 -1154
rect 1525 -1196 2482 -1192
rect 1332 -1218 1466 -1214
rect 1332 -1351 1336 -1218
rect 2478 -1223 2482 -1196
rect 384 -1381 1093 -1377
rect 2105 -1385 2515 -1381
rect 175 -1440 375 -1436
rect 175 -1616 179 -1440
rect 1432 -1653 2395 -1649
rect 86 -1844 122 -1840
rect -458 -1859 72 -1855
rect -1397 -2364 -471 -2360
rect -1397 -2706 -1393 -2364
rect -458 -2372 -454 -1859
rect -419 -1896 1357 -1892
rect -419 -2090 -415 -1896
rect 1432 -1895 1436 -1653
rect 2534 -1686 2538 -911
rect 3406 -1019 3410 -911
rect 2146 -1689 2538 -1686
rect 2146 -1690 2534 -1689
rect 2146 -2031 2150 -1690
rect -1388 -2376 -454 -2372
rect -1388 -2550 -1384 -2376
rect -105 -2578 -101 -2334
rect -586 -2582 -101 -2578
<< m3contact >>
rect -47 -57 -42 -52
rect -69 -111 -64 -106
rect 856 -265 861 -260
rect -122 -489 -117 -484
rect 619 -489 630 -483
rect -47 -500 -42 -495
rect -122 -883 -117 -878
rect 758 -490 763 -484
rect 931 -491 936 -486
rect 1372 -266 1378 -260
rect 1882 -266 1889 -260
rect 1341 -491 1346 -486
rect 1423 -492 1431 -487
rect 1649 -493 1654 -488
rect 780 -713 785 -708
rect 936 -1097 941 -1092
rect 959 -1097 964 -1091
rect 1671 -1236 1676 -1231
rect 2515 -1387 2521 -1379
rect 537 -1480 544 -1473
rect 1670 -1586 1676 -1581
rect 1578 -1620 1584 -1614
rect 936 -1726 941 -1721
rect 2867 -931 2873 -926
rect 2925 -1315 2930 -1310
rect -48 -1954 -43 -1949
rect 1614 -2007 1619 -2002
rect 2505 -1739 2510 -1734
rect 2609 -2123 2616 -2117
rect -834 -2415 -828 -2409
<< metal3 >>
rect -69 -177 -65 -111
rect -122 -181 -65 -177
rect -122 -484 -118 -181
rect -47 -252 -43 -57
rect -47 -256 1887 -252
rect -47 -476 -43 -256
rect -122 -878 -118 -489
rect -48 -495 -43 -476
rect -48 -500 -47 -495
rect -48 -1457 -44 -500
rect -834 -1461 -44 -1457
rect -834 -2409 -830 -1461
rect -48 -1949 -44 -1461
rect 537 -1473 541 -256
rect 630 -489 758 -485
rect 780 -708 784 -256
rect 856 -260 860 -256
rect 1372 -260 1376 -256
rect 936 -491 1341 -487
rect 959 -1091 963 -491
rect 1431 -492 1649 -488
rect 1671 -888 1675 -256
rect 1882 -260 1887 -256
rect 1671 -892 2872 -888
rect 936 -1615 940 -1097
rect 1671 -1231 1675 -892
rect 1671 -1581 1675 -1236
rect 936 -1619 1578 -1615
rect 936 -1721 940 -1619
rect 2505 -1734 2509 -892
rect 2868 -926 2872 -892
rect 2926 -1381 2930 -1315
rect 2521 -1385 2931 -1381
rect 1614 -2044 1618 -2007
rect 2610 -2044 2614 -1385
rect 1614 -2048 2614 -2044
rect 2610 -2117 2614 -2048
use and  and_0
timestamp 1638582313
transform 1 0 -6 0 1 -76
box 0 -34 56 24
use and  and_1
timestamp 1638582313
transform 1 0 120 0 1 -76
box 0 -34 56 24
use and  and_2
timestamp 1638582313
transform 1 0 246 0 1 -76
box 0 -34 56 24
use and  and_3
timestamp 1638582313
transform 1 0 372 0 1 -76
box 0 -34 56 24
use and  and_4
timestamp 1638582313
transform 1 0 498 0 1 -76
box 0 -34 56 24
use and  and_5
timestamp 1638582313
transform 1 0 624 0 1 -76
box 0 -34 56 24
use and  and_6
timestamp 1638582313
transform 1 0 750 0 1 -76
box 0 -34 56 24
use and  and_7
timestamp 1638582313
transform 1 0 876 0 1 -76
box 0 -34 56 24
use and  and_8
timestamp 1638582313
transform 1 0 1002 0 1 -76
box 0 -34 56 24
use and  and_9
timestamp 1638582313
transform 1 0 1128 0 1 -76
box 0 -34 56 24
use and  and_10
timestamp 1638582313
transform 1 0 1254 0 1 -76
box 0 -34 56 24
use and  and_11
timestamp 1638582313
transform 1 0 1380 0 1 -76
box 0 -34 56 24
use and  and_12
timestamp 1638582313
transform 1 0 1506 0 1 -76
box 0 -34 56 24
use and  and_13
timestamp 1638582313
transform 1 0 1632 0 1 -76
box 0 -34 56 24
use and  and_14
timestamp 1638582313
transform 1 0 1758 0 1 -76
box 0 -34 56 24
use and  and_15
timestamp 1638582313
transform 1 0 1884 0 1 -75
box 0 -34 56 24
use hadd  hadd_0
timestamp 1668432137
transform 1 0 846 0 1 -371
box -82 -121 126 112
use hadd  hadd_1
timestamp 1668432137
transform 1 0 1339 0 1 -372
box -82 -121 126 112
use hadd  hadd_2
timestamp 1668432137
transform 1 0 1850 0 1 -372
box -82 -121 126 112
use fadd  fadd_1
timestamp 1668441252
transform 1 0 -474 0 1 -727
box -71 -156 820 233
use fadd  fadd_0
timestamp 1668441252
transform 1 0 576 0 1 -940
box -71 -156 820 233
use fadd  fadd_5
timestamp 1668441252
transform 1 0 278 0 1 -1707
box -71 -156 820 233
use fadd  fadd_2
timestamp 1668441252
transform 1 0 1412 0 1 -1463
box -71 -156 820 233
use fadd  fadd_3
timestamp 1668441252
transform 1 0 2565 0 1 -1158
box -71 -156 820 233
use fadd  fadd_6
timestamp 1668441252
transform 1 0 -293 0 1 -2181
box -71 -156 820 233
use hadd  hadd_3
timestamp 1668432137
transform 1 0 1552 0 1 -1886
box -82 -121 126 112
use fadd  fadd_4
timestamp 1668441252
transform 1 0 2262 0 1 -1966
box -71 -156 820 233
use fadd  fadd_7
timestamp 1668441252
transform 1 0 -1279 0 1 -2641
box -71 -156 820 233
<< labels >>
rlabel metal1 -77 77 -69 81 4 A3
rlabel metal1 -77 66 -69 70 3 A2
rlabel metal1 -77 55 -69 59 3 A1
rlabel metal1 -77 44 -69 48 3 A0
rlabel metal1 -77 33 -69 37 3 B3
rlabel metal1 -77 22 -69 26 3 B2
rlabel metal1 -77 11 -69 15 3 B1
rlabel metal1 -77 0 -69 4 3 B0
rlabel metal1 61 -130 65 -124 1 and1
rlabel metal1 187 -130 191 -124 1 and2
rlabel metal1 313 -130 317 -124 1 and3
rlabel metal1 439 -130 443 -124 1 and4
rlabel metal1 565 -130 569 -124 1 and5
rlabel metal1 691 -130 695 -124 1 and6
rlabel metal1 817 -130 821 -124 1 and7
rlabel metal1 943 -130 947 -124 1 and8
rlabel metal1 1069 -130 1073 -124 1 and9
rlabel metal1 1195 -130 1199 -124 1 and10
rlabel metal1 1321 -130 1325 -124 1 and11
rlabel metal1 1447 -130 1451 -124 1 and12
rlabel metal1 1573 -130 1577 -124 1 and13
rlabel metal1 1699 -130 1703 -124 1 and14
rlabel metal1 1825 -130 1829 -124 1 and15
rlabel metal1 1951 -130 1955 -124 1 and16
rlabel metal1 -77 -110 -72 -106 3 gnd
rlabel metal1 -77 -56 -72 -52 3 vdd
rlabel metal1 4012 -2557 4016 -2548 7 P0
rlabel metal2 2026 -512 2030 -491 1 P1
rlabel metal1 3396 -1138 3405 -1134 1 P2
rlabel metal1 3095 -1946 3103 -1942 1 P3
rlabel metal1 1691 -1831 1699 -1827 1 P4
rlabel metal1 538 -2161 546 -2157 1 P5
rlabel metal1 -443 -2621 -436 -2617 1 P6
rlabel metal1 -448 -2507 -441 -2503 1 P7
<< end >>
